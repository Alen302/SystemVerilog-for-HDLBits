module zero (
    output var logic zero 
);
    
    assign zero = '0 ;
endmodule