module top_module (
    output var logic high
);

assign high = '1 ;
    
endmodule