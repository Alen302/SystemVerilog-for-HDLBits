module step_one (
    output var logic high
);

assign high = '1 ;
    
endmodule